`include "../../interfaces/PipelineInterface.svh"
`include "../core/utils/Opcodes.sv"
`include "../../interfaces/ControlSignals.svh"

module WB(
    input  logic clock,
    input  logic reset,
    input wire  mem_wb_bus_t mem_wb_bus_in,
    input wire  control_signals_t ctrl_signals_in
);

endmodule
