// Data structures for cache tag & data
parameter int TAGMSB = 19; // tag msb
parameter int TAGLSB = 6; // tag lsb


parameter int NUM_CACHE_BLOCKS = 4; // number of cache blocks
parameter int CACHE_BLOCK_SIZE = 128;  // cache block size (bytes)

parameter int NUM_MEM_BLOCKS = 1024; // number of memory blocks
parameter int MEM_BLOCK_SIZE = 128;  // memory block size (bytes)

parameter int NUM_PA_BITS = 10; // number of physical address bits


