parameter LW      = 7'b0000011;
parameter SW      = 7'b0100011;
parameter BEQ     = 7'b1100011;
parameter NOP_INST= 32'h00000013;
parameter ALUopR  = 7'b0110011; // R-type
parameter ALUopI  = 7'b0010011; // I-type
